module testbench();
	logic clk, reset;
	
	logic Tl, Tr, LA_expected, LB_expected, LC_expected, RA_expected, RB_expected, RC_expected;
	
	

endmodule