//// Модуль testbench тестирует другой модуль, испытываемое устройство(device under test).
// Он подает входные сигналы на ИУ и проверяет, соответствуют ли выходные сигналы ожидаемым значениям.
// Пользователь предоставляет шаблоны вводов и желаемых выводов, называемых testvectors (тестовые векторы).
module testbench();
	logic 		 clk, reset;
	// 'clk' & 'reset' - это частые имена для обозначения такта и сброса, но они не зарезервированы/
	logic 		 a, b, cin, s, cout, sexpected, coutexpected;
	// Эти переменные или сигналы представляют 3 ввода, 2 вывода, 2 ожидаемых вывода.
	logic [31:0] vectornum, errors;
	// '[31:0]' обозначает, что следующие сигналы,
	// "vectornum" и "errors" в этом случае являются 32-битными по длине (от 0 до 31 бит) в порядке от младшего к старшему 
	// (наименьший значащий бит по младшему адресу или [msb:lsb]). 
	// vectornum показывает количество применённых тестовых векторов.
	// errors показывает количество найденных ошибок.
	// Размер типа данных 'int' составляет 4 байта, таким образом 32 бита. 
	logic [4:0]  testvectors[10000:0];
	// Сверху вы можете видеть 5-битный двоичный массив, названный testvectors с индексом от 0 до 10000 
	//(testvectors[0],testvectors[1],testvectors[2],...,testvectors[10000]).
	// Другими словами, testvectors содержат 10001 элементов, каждый из которых - это 5-битное двоичное число. 
	// Количество битов представляет собой сумму количества входных и выходных битов
	// (к примеру. три 1-bit входа + два 1-битных выхода = один 5-битный testvector). 
	// В этом задании, мы будем использовать только 8 тестовых векторов (приведен ниже .tv),
	// однако не ничего страшного в том, чтобы установить массив для использования большего количества, 
	// так что мы сможем спокойно добавить тестовые векторы позже.

//// Инстанцируем испытываемое устройство (ИУ/DUT).
// Входы: a, b, cin. выходы: s, cout.
fulladder dut(a, b, cin, s, cout);

//// Тактовый генератор синхросигнала.
always
// Оператор 'always' заставляет утверждения в блоке постоянно переоцениваться.
	begin
      	//// Создать такт с периодом 10 единиц времени. 
		// Назначить сигнал clk HIGH(1) на 5 единиц, LOW(0) на 5 единиц 
		clk=1; #5; 
		clk=0; #5;
	end

//// Начало теста. 
initial
// 'initial' используется только в симуляции (несинтезируемое подмножество).
	begin
		//// Загрузить векторы, хранящиеся как нули и единицы (в двоичном формате) в .tv-файле.
		$readmemb("fulladder.tv", testvectors);
		// $readmemb читает двоичный формат, $readmemh читает шестнадцатеричный формат.

		// Инициализировать количество применённых векторов и количество обнаруженных ошибок.
		vectornum=0; 
		errors=0;
		// Оба сигнала инициализированы нулями в начале.

		//// Сброс импульса на 22 единицы времени (2,2 цикла), поэтому сигнал reset падает после фронта синхросигнала.
		reset=1; #22;
     	reset=0;
		// Сигнал становится HIGH(1) на 22 единицы времени, затем остается LOW(0) до конца теста.
	end

//// Применяйте тестовые векторы по нарастающему фронту сигнала clk.
always @(posedge clk)
	//  Обратите внимание, что этот оператор 'always' имеет список чувствительности,
	// который контролирует, когда все утверждения в блоке начнут оцениваться. 
	// '@(posedge clk)' означает по положительному или нарастающему фронту тактового cигнала. 
	begin
		//// Применяйте тестовые векторы через 1 единицу времени после нарастающего фронта тактового сигнала,
		// чтобы избежать изменения данных одновременно с тактовым сигналом.
		#1;
		//// Разбейте текущий 5-битный тестовый вектор на 3 входа и 2 ожидаемых выхода.
 		{a,b,cin, coutexpected,sexpected} = testvectors[vectornum];
	end

//// Проверка результатов по спадающему фронту сигнала clk.
always @(negedge clk)
// Эта строка кода позволяет программе выполнить следующие утверждения
// в блоке по отрицательному фронту тактового сигнала.
	//// Ничего не делает во время сброса. В противном случае проверяете результат.
	if (~reset) begin
			//// Находит ошибки, проверяя если выводы из ИУ совпадают с ожиданиями.
			if (s !== sexpected || cout !== coutexpected) begin
			// Если обнаружена ошибка, выводит все 3 входа, 2 выхода, 2 ожидаемых выхода.
				$display("Error: inputs = %b", {a, b, cin});
				// '$display' выводит любое утверждение внутри кавычек в окно симулятора.
				// %b, %d и %h указывают значения в двоичном, десятичном и шестнадцатеричном форматах.
				// {a, b, cin} создают вектор, содержащий три сигнала.
				$display(" outputs = %b %b (%b %b expected)", s, cout, sexpected, coutexpected);
				//// Увеличивает количество errors.
				errors = errors + 1;
			end
			//// Увеличиваем количество векторов.
			vectornum = vectornum + 1;
			//// Когда вектор теста становится равным 'x', это означает, что все векторы,
            // которые были первоначально загружены, были обработаны, и таким образом тест завершен.
			if (testvectors[vectornum] === 5'bx) begin
			// '==='&'!==' может сравнивать неизвестные и плавающие значения (X&Z),
			// в отличие от. '=='&'!=', который может сравнивать только 0 и 1.
			// 5'bx - 5-битное двоичное число x или xxxxx.
			// Если текущий тестовый вектор равен xxxxx, сообщает количество векторов и обнаруженных ошибок.
				$display("%d tests completed with %d errors", vectornum, errors);
				// Затем остановите симуляцию.
			$stop;
		end
	end

// Резюмируя, новые входы подаются по положительному фронту тактового сигнала
// и выходы проверяются на соответствие ожидаемым выходам на отрицательном тактовом сигнале. 
// Об ошибках сообщается одновременно. 
// Процесс повторяется до тех пор, пока в массивах testvectors не останется допустимых тестовых векторов. 
// В конце симулирования модуль выводит общее количество примененных тестовых векторов и общее количество обнаруженных ошибок. 
endmodule